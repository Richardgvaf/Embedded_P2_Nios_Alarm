// prueba1_tb.v

// Generated using ACDS version 19.1 670

`timescale 1 ps / 1 ps
module prueba1_tb (
	);

	wire        prueba1_inst_clk_bfm_clk_clk;                                       // prueba1_inst_clk_bfm:clk -> [prueba1_inst:clk_clk, prueba1_inst_reset_bfm:clk]
	wire  [2:0] prueba1_inst_button_input_1_external_connection_bfm_conduit_export; // prueba1_inst_button_input_1_external_connection_bfm:sig_export -> prueba1_inst:button_input_1_external_connection_export
	wire  [7:0] prueba1_inst_led_output_5_external_connection_export;               // prueba1_inst:led_output_5_external_connection_export -> prueba1_inst_led_output_5_external_connection_bfm:sig_export
	wire  [7:0] prueba1_inst_regs_export;                                           // prueba1_inst:regs_export -> prueba1_inst_regs_bfm:sig_export
	wire  [7:0] prueba1_inst_ss_output_1_external_conection_export;                 // prueba1_inst:ss_output_1_external_conection_export -> prueba1_inst_ss_output_1_external_conection_bfm:sig_export
	wire  [7:0] prueba1_inst_ss_output_2_external_connection_export;                // prueba1_inst:ss_output_2_external_connection_export -> prueba1_inst_ss_output_2_external_connection_bfm:sig_export
	wire  [7:0] prueba1_inst_ss_output_3_external_connection_export;                // prueba1_inst:ss_output_3_external_connection_export -> prueba1_inst_ss_output_3_external_connection_bfm:sig_export
	wire  [7:0] prueba1_inst_ss_output_4_external_connection_export;                // prueba1_inst:ss_output_4_external_connection_export -> prueba1_inst_ss_output_4_external_connection_bfm:sig_export
	wire  [2:0] prueba1_inst_switch_input_2_external_connection_bfm_conduit_export; // prueba1_inst_switch_input_2_external_connection_bfm:sig_export -> prueba1_inst:switch_input_2_external_connection_export
	wire        prueba1_inst_reset_bfm_reset_reset;                                 // prueba1_inst_reset_bfm:reset -> prueba1_inst:reset_reset_n

	prueba1 prueba1_inst (
		.button_input_1_external_connection_export (prueba1_inst_button_input_1_external_connection_bfm_conduit_export), // button_input_1_external_connection.export
		.clk_clk                                   (prueba1_inst_clk_bfm_clk_clk),                                       //                                clk.clk
		.led_output_5_external_connection_export   (prueba1_inst_led_output_5_external_connection_export),               //   led_output_5_external_connection.export
		.regs_export                               (prueba1_inst_regs_export),                                           //                               regs.export
		.reset_reset_n                             (prueba1_inst_reset_bfm_reset_reset),                                 //                              reset.reset_n
		.ss_output_1_external_conection_export     (prueba1_inst_ss_output_1_external_conection_export),                 //     ss_output_1_external_conection.export
		.ss_output_2_external_connection_export    (prueba1_inst_ss_output_2_external_connection_export),                //    ss_output_2_external_connection.export
		.ss_output_3_external_connection_export    (prueba1_inst_ss_output_3_external_connection_export),                //    ss_output_3_external_connection.export
		.ss_output_4_external_connection_export    (prueba1_inst_ss_output_4_external_connection_export),                //    ss_output_4_external_connection.export
		.switch_input_2_external_connection_export (prueba1_inst_switch_input_2_external_connection_bfm_conduit_export)  // switch_input_2_external_connection.export
	);

	altera_conduit_bfm prueba1_inst_button_input_1_external_connection_bfm (
		.sig_export (prueba1_inst_button_input_1_external_connection_bfm_conduit_export)  // conduit.export
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) prueba1_inst_clk_bfm (
		.clk (prueba1_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_conduit_bfm_0002 prueba1_inst_led_output_5_external_connection_bfm (
		.sig_export (prueba1_inst_led_output_5_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0002 prueba1_inst_regs_bfm (
		.sig_export (prueba1_inst_regs_export)  // conduit.export
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) prueba1_inst_reset_bfm (
		.reset (prueba1_inst_reset_bfm_reset_reset), // reset.reset_n
		.clk   (prueba1_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_conduit_bfm_0002 prueba1_inst_ss_output_1_external_conection_bfm (
		.sig_export (prueba1_inst_ss_output_1_external_conection_export)  // conduit.export
	);

	altera_conduit_bfm_0002 prueba1_inst_ss_output_2_external_connection_bfm (
		.sig_export (prueba1_inst_ss_output_2_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0002 prueba1_inst_ss_output_3_external_connection_bfm (
		.sig_export (prueba1_inst_ss_output_3_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm_0002 prueba1_inst_ss_output_4_external_connection_bfm (
		.sig_export (prueba1_inst_ss_output_4_external_connection_export)  // conduit.export
	);

	altera_conduit_bfm prueba1_inst_switch_input_2_external_connection_bfm (
		.sig_export (prueba1_inst_switch_input_2_external_connection_bfm_conduit_export)  // conduit.export
	);

endmodule
